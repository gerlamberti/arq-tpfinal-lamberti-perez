`timescale 1ns/1ps

module IF_EX #()();




endmodule