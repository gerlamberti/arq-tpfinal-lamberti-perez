
// Opcodes
`define RTYPE_OPCODE 6'b000000
`define ADDI_OPCODE 6'b001000




// Function codes for R-type instructions
`define ADD_FCODE 6'b100000
`define ADDU_FCODE 6'b100001
`define AND_FCODE 6'b100100
`define JALR_FCODE 6'b001001
`define NOR_FCODE 6'b100111
`define OR_FCODE 6'b100101
`define SLL_FCODE 6'b000000
`define SLLV_FCODE 6'b000100
`define SLT_FCODE 6'b101010
`define SRA_FCODE 6'b000011
`define SRAV_FCODE 6'b000111
`define SRL_FCODE 6'b000010
`define SRLV_FCODE 6'b000110
`define SUB_FCODE 6'b100010
`define SUBU_FCODE 6'b100011
`define XOR_FCODE 6'b100110

