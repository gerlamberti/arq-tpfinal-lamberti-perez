// Word Size params
`define COMPLETE_WORD   3'b100
`define HALF_WORD       3'b010
`define BYTE_WORD       3'b001