`timescale 1ns/1ps

module register_file #()();




endmodule