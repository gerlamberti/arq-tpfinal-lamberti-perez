// Extensions Mode
`define SIGNED_EXTENSION_MODE 2'b00
`define UNSIGNED_EXTENSION_MODE 2'b01
`define SHIFT16L_EXTENSION_MODE 2'b10

// ALU SRC
`define RT_ALU_SRC 1'b0
`define INMEDIATE_ALU_SRC 1'b1
