`timescale 1ns/1ps

module ID #()();




endmodule